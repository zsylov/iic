library verilog;
use verilog.vl_types.all;
entity IIC_demo_vlg_tst is
end IIC_demo_vlg_tst;
